`ifdef RTL
    `define CYCLE_TIME 6.0
`endif
`ifdef GATE
    `define CYCLE_TIME 6.0
`endif


`define PATNUM 10

module PATTERN(
    // Output signals
    clk,
 rst_n,
 in_valid,
    in_data, 
 in_mode,
    // Input signals
    out_valid, 
 out_data
);

// ========================================
// Input & Output
// ========================================
output reg clk, rst_n, in_valid;
output reg [8:0] in_mode;
output reg [14:0] in_data;

input out_valid;
input [206:0] out_data;

//================================================================
// clock
//================================================================
real CYCLE = `CYCLE_TIME;
always #(CYCLE/2.0) clk = ~clk;
initial clk = 0;

integer PATNUM = `PATNUM;
integer patcount;
integer latency, total_latency;
localparam [8:0] in_mode_array [0:2] = {9'b010101000, 9'b100001100, 9'b011001100};
integer mode_idx;
integer file;

reg signed[206:0] golden_outdata;


reg signed [10:0] golden_in_data[0:3][0:3];
reg [14:0] in_data_temp[0:3][0:3];
reg signed [22:0] out_temp_two_by_two[0:8];
reg signed [50:0] out_temp_three_by_three[0:3];
reg signed [206:0] out_temp_four_by_four;
reg signed [206:0] si_out_data;
reg [8:0] in_mode_temp;
reg [8:0] in_mode_flip;
reg signed [22:0] your_out_2 [0:8];
reg signed [50:0] your_out_3 [0:3];


reg [4:0] golden_in_mode;
reg [4:0] error_bit;
reg [3:0] flip_bit;



/* Check for invalid overlap */
always @(*) begin
    if (in_valid && out_valid) begin
        display_fail;
        $display("************************************************************");  
        $display("                          FAIL!                           ");    
        $display("*  The out_valid signal cannot overlap with in_valid.   *");
        $display("************************************************************");
        $finish;            
    end    
end



initial begin

    reset_task;
    file = $fopen("../00_TESTBED/debug.txt", "w");
 for( patcount = 0; patcount < PATNUM; patcount++) begin 
        repeat($urandom_range(2,4)) @(negedge clk); 
        input_task;
        write_input_to_file;
        wait_out_valid_task;
  check_ans;
        $display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32mExecution Cycle: %3d, \033[0;33m", patcount + 1, latency);
  
 end
 display_pass;
    repeat(3) @(negedge clk);
    $finish;
end





task reset_task; begin 
    rst_n = 1'b1;
    in_valid = 1'b0;
    in_data = 15'bx;
    in_mode = 9'bx;
    total_latency = 0;

    force clk = 0;

    // Apply reset
    #CYCLE; rst_n = 1'b0; 
    #CYCLE; rst_n = 1'b1;
    
    // Check initial conditions
    if (out_valid !== 1'b0 || out_data !== 'b0) begin
        display_fail;
        $display("************************************************************");  
        $display("                          FAIL!                           ");    
        $display("*  Output signals should be 0 after initial RESET at %8t *", $time);
        $display("************************************************************");
        repeat (2) #CYCLE;
        $finish;
    end
    #CYCLE; release clk;
end endtask



task input_task; begin
    integer i,j;
    in_valid = 1'b1;
    for(i = 0; i < 16; i = i + 1) begin
        in_data = $urandom_range(0, 32767);   // 15-bit random data
        in_data_temp[i / 4][i % 4] = in_data;
        if(i == 0)begin
            mode_idx = $urandom_range(0, 2);
            in_mode_flip = in_mode_array[mode_idx];
            $display("correct: %b",{in_mode_flip[6],in_mode_flip[4],in_mode_flip[3],in_mode_flip[2],in_mode_flip[0]});
            flip_bit = $urandom_range(0, 10);
            if(flip_bit < 9)begin
                in_mode_flip[5 + 4 - flip_bit] = ~in_mode_flip[5 + 4 - flip_bit];
            end
            in_mode = in_mode_flip;
            in_mode_temp = in_mode_flip;
            //decode mode here!
            error_bit = 0;
            for(j = 0; j < 5 + 4; j = j + 1) begin
                if(in_mode_flip[5 + 4 - j - 1] === 1'b1)begin
                    error_bit = error_bit ^ (j + 1);
                end
            end
            in_mode_flip[5 + 4 - error_bit] = ~in_mode_flip[5 + 4 - error_bit];
            golden_in_mode = {in_mode_flip[6],in_mode_flip[4],in_mode_flip[3],in_mode_flip[2],in_mode_flip[0]};

        end
        else begin
            in_mode = 'bx;
        end
        @(negedge clk);
    end
    in_data_decode;
    in_data = 15'bx;
    in_mode = 9'bx;
    in_valid = 1'b0;
   
    
end endtask


task wait_out_valid_task; begin
    latency = 0;
    while (out_valid !== 1'b1) begin
        latency = latency + 1;
        if (latency == 1000) begin
            display_fail;
            $display("********************************************************");     
            $display("                          FAIL!                           ");
            $display("*  The execution latency exceeded 1000 cycles at %8t   *", $time);
            $display("********************************************************");
            repeat (2) @(negedge clk);
            $finish;
        end
        @(negedge clk);
    end
    total_latency = total_latency + latency;
end endtask



task check_ans; begin
    si_out_data = out_data;
    calculate_golden_outdata;
    write_output_to_file;
    

    if (out_data !== golden_outdata) begin
        if (golden_in_mode == 5'b00100) begin
            $display ("                          matrix size is 2*2                  ");
            $display ("            determinant should be : %d\t%d\t%d           ", out_temp_two_by_two[0], out_temp_two_by_two[1], out_temp_two_by_two[2]);
            $display ("                                    %d\t%d\t%d           ", out_temp_two_by_two[3], out_temp_two_by_two[4], out_temp_two_by_two[5]);
            $display ("                                    %d\t%d\t%d           ", out_temp_two_by_two[6], out_temp_two_by_two[7], out_temp_two_by_two[8]);
            $display ("            your answer is        : %d\t%d\t%d           ",  out_data[206:184], out_data[183:161], out_data[160:138]);
            $display ("                                    %d\t%d\t%d           ", out_data[137:115], out_data[114:92], out_data[91:69]);
            $display ("                                    %d\t%d\t%d           ", out_data[68:46], out_data[45:23], out_data[22:0]);
        end
        else if (golden_in_mode == 5'b00110) begin
            $display ("                          matrix size is 3*3                  ");
            $display ("            determinant should be : %d\t%d           ", out_temp_three_by_three[0], out_temp_three_by_three[1]);
            $display ("                                    %d\t%d           ", out_temp_three_by_three[2], out_temp_three_by_three[3]);
            $display ("            your answer is        : %d\t%d           ", out_data[203:153], out_data[152:102]);
            $display ("                                    %d\t%d           ", out_data[101:51], out_data[50:0]);
        end 
        else begin
            $display ("                          matrix size is 4*4                  ");
            $display ("            determinant should be : %d           ", out_temp_four_by_four);
            $display ("            your answer is        : %d           ", si_out_data);
        end
        repeat (9) @(negedge clk);
        $finish;
    end
    

    @(negedge clk);
        
    // Check if the number of outputs matches the expected count
    if(out_valid === 1'b1) begin
        display_fail;
        $display("************************************************************");  
        $display("                          FAIL!                              ");
        $display("                Expected one valid output                    ");
        $display("************************************************************");
        repeat(9) @(negedge clk);
        $finish;
    end
end endtask



// task mode_decode;begin
//     integer i;
//     for(integer i = 0; i < 5 + 4; i = i + 1) begin
//         error_bit = 0;
//         if(in_mode_temp[5 + 4 - i - 1] === 1'b1)begin
//             error_bit = error_bit ^ (i + 1);
//         end
//     end
//     $display("%d",error_bit);
//     $display("func in: %b",in_mode_temp[i]);
//     in_mode_temp[5 + 4 - error_bit] = ~in_mode_temp[5 + 4 - error_bit];
//     golden_in_mode = {in_mode_temp[6],in_mode_temp[4],in_mode_temp[3],in_mode_temp[2],in_mode_temp[0]};
//     $display("func out :%b",golden_in_mode[i]);
// end endtask





task in_data_decode;begin
    for(integer i = 0; i < 4 ; i = i + 1)begin
        for(integer j = 0; j < 4 ; j = j + 1)begin
            error_bit = 0;
            for(integer k = 0; k < 11 + 4; k = k + 1) begin
                if(in_data_temp[i][j][11 + 4 - k - 1] === 1'b1)begin
                    error_bit = error_bit ^ (k + 1);
                end
            end
            // $display("%d",error_bit);
            // $display("in: %b",in_data_temp[i][j]);
            in_data_temp[i][j][11 + 4 - error_bit] = ~in_data_temp[i][j][11 + 4 - error_bit];

            golden_in_data[i][j] = {in_data_temp[i][j][12],in_data_temp[i][j][10],in_data_temp[i][j][9],in_data_temp[i][j][8],
                in_data_temp[i][j][6],in_data_temp[i][j][5],in_data_temp[i][j][4],in_data_temp[i][j][3],in_data_temp[i][j][2],
                in_data_temp[i][j][1],in_data_temp[i][j][0]};
            // $display("out :%b",golden_in_data[i][j]);
        end 
    end
end endtask

task calculate_golden_outdata;begin
    

    out_temp_two_by_two[0] = golden_in_data[0][0] * golden_in_data[1][1] - golden_in_data[0][1] * golden_in_data[1][0];
    out_temp_two_by_two[1] = golden_in_data[0][1] * golden_in_data[1][2] - golden_in_data[0][2] * golden_in_data[1][1];
    out_temp_two_by_two[2] = golden_in_data[0][2] * golden_in_data[1][3] - golden_in_data[0][3] * golden_in_data[1][2];
    out_temp_two_by_two[3] = golden_in_data[1][0] * golden_in_data[2][1] - golden_in_data[1][1] * golden_in_data[2][0];
    out_temp_two_by_two[4] = golden_in_data[1][1] * golden_in_data[2][2] - golden_in_data[1][2] * golden_in_data[2][1];
    out_temp_two_by_two[5] = golden_in_data[1][2] * golden_in_data[2][3] - golden_in_data[1][3] * golden_in_data[2][2];
    out_temp_two_by_two[6] = golden_in_data[2][0] * golden_in_data[3][1] - golden_in_data[2][1] * golden_in_data[3][0];
    out_temp_two_by_two[7] = golden_in_data[2][1] * golden_in_data[3][2] - golden_in_data[2][2] * golden_in_data[3][1];
    out_temp_two_by_two[8] = golden_in_data[2][2] * golden_in_data[3][3] - golden_in_data[2][3] * golden_in_data[3][2];

    out_temp_three_by_three[0] = golden_in_data[0][0] * golden_in_data[1][1] * golden_in_data[2][2] +
                                golden_in_data[0][1] * golden_in_data[1][2] * golden_in_data[2][0] +
                                golden_in_data[0][2] * golden_in_data[1][0] * golden_in_data[2][1] -
                                golden_in_data[0][2] * golden_in_data[1][1] * golden_in_data[2][0] -
                                golden_in_data[1][2] * golden_in_data[2][1] * golden_in_data[0][0] -
                                golden_in_data[0][1] * golden_in_data[1][0] * golden_in_data[2][2];
    
    out_temp_three_by_three[1] = golden_in_data[0][1] * golden_in_data[1][2] * golden_in_data[2][3] +
                                golden_in_data[0][2] * golden_in_data[1][3] * golden_in_data[2][1] +
                                golden_in_data[0][3] * golden_in_data[1][1] * golden_in_data[2][2] -
                                golden_in_data[0][3] * golden_in_data[1][2] * golden_in_data[2][1] -
                                golden_in_data[1][3] * golden_in_data[2][2] * golden_in_data[0][1] -
                                golden_in_data[0][2] * golden_in_data[1][1] * golden_in_data[2][3];
    
    out_temp_three_by_three[2] = golden_in_data[1][0] * golden_in_data[2][1] * golden_in_data[3][2] +
                                golden_in_data[1][1] * golden_in_data[2][2] * golden_in_data[3][0] +
                                golden_in_data[1][2] * golden_in_data[2][0] * golden_in_data[3][1] -
                                golden_in_data[1][2] * golden_in_data[2][1] * golden_in_data[3][0] -
                                golden_in_data[2][2] * golden_in_data[3][1] * golden_in_data[1][0] -
                                golden_in_data[1][1] * golden_in_data[2][0] * golden_in_data[3][2];

    out_temp_three_by_three[3] = golden_in_data[1][1] * golden_in_data[2][2] * golden_in_data[3][3] +
                                golden_in_data[1][2] * golden_in_data[2][3] * golden_in_data[3][1] +
                                golden_in_data[1][3] * golden_in_data[2][1] * golden_in_data[3][2] -
                                golden_in_data[1][3] * golden_in_data[2][2] * golden_in_data[3][1] -
                                golden_in_data[2][3] * golden_in_data[3][2] * golden_in_data[1][1] -
                                golden_in_data[1][2] * golden_in_data[2][1] * golden_in_data[3][3];
    
out_temp_four_by_four = golden_in_data[0][0] * (
                golden_in_data[1][1] * golden_in_data[2][2] * golden_in_data[3][3] +
                golden_in_data[1][2] * golden_in_data[2][3] * golden_in_data[3][1] +
                golden_in_data[1][3] * golden_in_data[2][1] * golden_in_data[3][2] -
                golden_in_data[1][3] * golden_in_data[2][2] * golden_in_data[3][1] -
                golden_in_data[1][2] * golden_in_data[2][1] * golden_in_data[3][3] -
                golden_in_data[1][1] * golden_in_data[2][3] * golden_in_data[3][2])
            - golden_in_data[0][1] * (
                golden_in_data[1][0] * golden_in_data[2][2] * golden_in_data[3][3] +
                golden_in_data[1][2] * golden_in_data[2][3] * golden_in_data[3][0] +
                golden_in_data[1][3] * golden_in_data[2][0] * golden_in_data[3][2] -
                golden_in_data[1][3] * golden_in_data[2][2] * golden_in_data[3][0] -
                golden_in_data[1][2] * golden_in_data[2][0] * golden_in_data[3][3] -
                golden_in_data[1][0] * golden_in_data[2][3] * golden_in_data[3][2])
            + golden_in_data[0][2] * (
                golden_in_data[1][0] * golden_in_data[2][1] * golden_in_data[3][3] +
                golden_in_data[1][1] * golden_in_data[2][3] * golden_in_data[3][0] +
                golden_in_data[1][3] * golden_in_data[2][0] * golden_in_data[3][1] -
                golden_in_data[1][3] * golden_in_data[2][1] * golden_in_data[3][0] -
                golden_in_data[1][1] * golden_in_data[2][0] * golden_in_data[3][3] -
                golden_in_data[1][0] * golden_in_data[2][3] * golden_in_data[3][1])
             - golden_in_data[0][3] * (
                golden_in_data[1][0] * golden_in_data[2][1] * golden_in_data[3][2] +
                golden_in_data[1][1] * golden_in_data[2][2] * golden_in_data[3][0] +
                golden_in_data[1][2] * golden_in_data[2][0] * golden_in_data[3][1] -
                golden_in_data[1][2] * golden_in_data[2][1] * golden_in_data[3][0] -
                golden_in_data[1][1] * golden_in_data[2][0] * golden_in_data[3][2] -
                golden_in_data[1][0] * golden_in_data[2][2] * golden_in_data[3][1]);

                                
    

    if(golden_in_mode == 5'b00100)begin
        golden_outdata = {out_temp_two_by_two[0],out_temp_two_by_two[1],out_temp_two_by_two[2],out_temp_two_by_two[3],out_temp_two_by_two[4],out_temp_two_by_two[5],out_temp_two_by_two[6],out_temp_two_by_two[7],out_temp_two_by_two[8]};
    end
    else if(golden_in_mode == 5'b00110)begin
        
        golden_outdata = {3'b000, out_temp_three_by_three[0],out_temp_three_by_three[1],out_temp_three_by_three[2],out_temp_three_by_three[3]};
    end
    else if(golden_in_mode == 5'b10110)begin
        golden_outdata = out_temp_four_by_four;
    end
    
end endtask


task write_input_to_file; begin
    $fwrite(file, "===========  PATTERN NO.%4d  ====\n", patcount);
    $fwrite(file, "===========  in_mode = %5b  =====\n",golden_in_mode);
    $fwrite(file, "===========  in_data  ===========\n");
    for(integer i = 0; i < 4; i = i + 1) begin
        for(integer j = 0; j < 4; j = j + 1) begin
            $fwrite(file, "%7d ", golden_in_data[i][j]);
        end
        $fwrite(file, "\n");
    end
    $fwrite(file, "===========   out_data   ==========\n");

end endtask

task write_output_to_file; begin
    $fwrite(file, "===========  2 * 2   =========\n");
    for(integer i = 0; i < 9; i = i + 1) begin
        $fwrite(file, "%10d ", out_temp_two_by_two[i]);
        if(i % 3 == 2)begin
            $fwrite(file, "\n");
        end
    end
    $fwrite(file, "===========  3 * 3   ========\n");
    for(integer i = 0; i < 4; i = i + 1) begin
        $fwrite(file, "%15d", out_temp_three_by_three[i]);
        if(i % 2 == 1)begin
            $fwrite(file, "\n");
        end
    end
    $fwrite(file, "===========  4 * 4   =========\n");
    $fwrite(file, "%20d\n", out_temp_four_by_four);

    $fwrite(file, "==========  golden out_data  ========\n");
    $fwrite(file, "%20d\n\n\n\n\n", golden_outdata);
end endtask







task display_fail; begin
    $display("\n");
    $display("\n");
    $display("\033[0;37m....................................................................................................\033[0m");
    $display("\033[0;37m.......................................................................,:+++:.......................\033[0m");
    $display("\033[0;37m....................................................,:+*\033[0m\033[0;32m******\033[0m\033[0;37m+;,....:*\033[0m\033[0;30m%%%%?%%S\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m*:....................\033[0m");
    $display("\033[0;37m................................................,:*\033[0m\033[0;30m?%%%%%%%%\033[0m\033[0;32m????\033[0m\033[0;30m?%%%%%%%%\033[0m\033[0;32m*\033[0m\033[0;37m:.;.\033[0m\033[0;30m%%\033[0m\033[0;32m?\033[0m\033[0;30m%%SS%%%%SSS%%\033[0m\033[0;37m:..................\033[0m");
    $display("\033[0;37m..............................................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m?????\033[0m\033[0;30m%%SSSSSSSSSSS\033[0m\033[0;37m.\033[0m\033[0;30m%%%%SSSSSS%%%%%%S\033[0m\033[0;37m.*,................\033[0m");
    $display("\033[0;37m...........................................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m??????\033[0m\033[0;30mSS%%%%%%%%SSSSS#\033[0m\033[0;37m..\033[0m\033[0;30mSSSSS%%\033[0m\033[0;32m???????\033[0m\033[0;30m%%SS\033[0m\033[0;37m;...............\033[0m");
    $display("\033[0;37m........................................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m???????\033[0m\033[0;30m%%S%%?%%SS%%%%???%%%%%%\033[0m\033[0;37m..\033[0m\033[0;30mSS%%\033[0m\033[0;32m??\033[0m\033[0;30m%%%%%%%%?\033[0m\033[0;32m*\033[0m\033[0;37m***\033[0m\033[0;30m?S\033[0m\033[0;37m*..............\033[0m");
    $display("\033[0;37m....................................,:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m????????\033[0m\033[0;30m%%SS?%%S%%\033[0m\033[0;32m???????????\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;30m%%?%%?\033[0m\033[0;37m+:,.,;+;,.,+\033[0m\033[0;30m?\033[0m\033[0;37m,............\033[0m");
    $display("\033[0;37m.................................,;*\033[0m\033[0;30m?%%?\033[0m\033[0;32m???????????\033[0m\033[0;30m%%\033[0m\033[0;32m?\033[0m\033[0;30m%%S%%\033[0m\033[0;32m????????\033[0m\033[0;30m?%%%%%%%%%%S\033[0m\033[0;37m.+:....+.....+..*\033[0m\033[0;30m*\033[0m\033[0;37m............\033[0m");
    $display("\033[0;37m..............................,;\033[0m\033[0;32m*\033[0m\033[0;30m%%%%?\033[0m\033[0;32m???????????????\033[0m\033[0;30mSS\033[0m\033[0;32m???????\033[0m\033[0;30m%%%%?\033[0m\033[0;32m*\033[0m\033[0;37m*+++++\033[0m\033[0;30mS\033[0m\033[0;37m,....:.......:..\033[0m\033[0;30mS\033[0m\033[0;37m:...........\033[0m");
    $display("\033[0;37m...........................:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m??????????????????\033[0m\033[0;30m%%S\033[0m\033[0;32m????\033[0m\033[0;30m%%%%%%?\033[0m\033[0;37m+;::,.....\033[0m\033[0;30mS\033[0m\033[0;37m;....*....;\033[0m\033[0;30m?\033[0m\033[0;37m.\033[0m\033[0;30m?\033[0m\033[0;37m,+.+...........\033[0m");
    $display("\033[0;37m.......................,:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m?????????????????????\033[0m\033[0;30mSS%%%%%%%%\033[0m\033[0;32m*\033[0m\033[0;37m;,,\033[0m\033[0;30m?\033[0m\033[0;37m....*.....\033[0m\033[0;30mS\033[0m\033[0;37m:,..\033[0m\033[0;30m?\033[0m\033[0;37m....;\033[0m\033[0;30m?\033[0m\033[0;37m..\033[0m\033[0;30m%%%%%%\033[0m\033[0;37m;...........\033[0m");
    $display("\033[0;37m....................,:+\033[0m\033[0;30m?%%%%\033[0m\033[0;32m???????????????????????\033[0m\033[0;30m%%%%S\033[0m\033[0;37m;:,,..:.......+..;.\033[0m\033[0;30m#SS%%?S\033[0m\033[0;37m.....\033[0m\033[0;30mS%%SS\033[0m\033[0;37m.*............\033[0m");
    $display("\033[0;37m..................,+\033[0m\033[0;30m?%%?\033[0m\033[0;32m??????????????????????????\033[0m\033[0;30m%%S?%%\033[0m\033[0;37m;...,....+\033[0m\033[0;30m%%\033[0m\033[0;37m..\033[0m\033[0;30m%%\033[0m\033[0;37m.+..\033[0m\033[0;30m%%\033[0m\033[0;32m*?\033[0m\033[0;30mSSSSSS%%SS\033[0m\033[0;37m....\033[0m\033[0;30m?\033[0m\033[0;37m,...........\033[0m");
    $display("\033[0;37m................:*\033[0m\033[0;30m??\033[0m\033[0;32m????????????????????????\033[0m\033[0;30m#?\033[0m\033[0;32m????\033[0m\033[0;30m#%%\033[0m\033[0;32m?\033[0m\033[0;30mS%%\033[0m\033[0;37m*:\033[0m\033[0;30m?\033[0m\033[0;37m...\033[0m\033[0;35m*\033[0m\033[0;37m,\033[0m\033[0;30m?\033[0m\033[0;37m...\033[0m\033[0;30mSS?%%\033[0m\033[0;37m..\033[0m\033[0;30m%%?\033[0m\033[0;32m?????\033[0m\033[0;30m%%SS#S%%\033[0m\033[0;32m?\033[0m\033[0;30m%%\033[0m\033[0;33m*\033[0m\033[0;37m...........\033[0m");
    $display("\033[0;37m..............,*\033[0m\033[0;30m%%\033[0m\033[0;32m???????????????????????????\033[0m\033[0;37m..\033[0m\033[0;30m%%\033[0m\033[0;32m????\033[0m\033[0;30m#S\033[0m\033[0;32m??\033[0m\033[0;30m%%S#\033[0m\033[0;37m...\033[0m\033[0;30mSS\033[0m\033[0;37m.\033[0m\033[0;30m#SS%%\033[0m\033[0;32m????\033[0m\033[0;30m%%\033[0m\033[0;37m...\033[0m\033[0;30mSSSSS%%?\033[0m\033[0;32m?????\033[0m\033[0;30m%%\033[0m\033[0;37m,..........\033[0m");
    $display("\033[0;37m.............+\033[0m\033[0;30m%%?\033[0m\033[0;32m?????????????????????????????\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;30m#%%%%\033[0m\033[0;32m??\033[0m\033[0;30m%%SSSSSS%%SSS%%%%\033[0m\033[0;32m?????????\033[0m\033[0;30m%%\033[0m\033[0;37m..\033[0m\033[0;30mS%%\033[0m\033[0;32m?????????\033[0m\033[0;30m%%\033[0m\033[0;37m,..........\033[0m");
    $display("\033[0;37m............*\033[0m\033[0;30mS\033[0m\033[0;32m??????\033[0m\033[0;30m%%%%%%\033[0m\033[0;32m????\033[0m\033[0;30m%%%%%%%%%%%%%%%%%%%%%%%%?\033[0m\033[0;32m???????\033[0m\033[0;30m?%%SSSSSSS##S%%%%?\033[0m\033[0;32m??????????????\033[0m\033[0;30mS%%\033[0m\033[0;32m???????\033[0m\033[0;30m?%%%%\033[0m\033[0;37m+...........\033[0m");
    $display("\033[0;37m...........:\033[0m\033[0;30mS\033[0m\033[0;32m??????\033[0m\033[0;30m%%%%\033[0m\033[0;32m???\033[0m\033[0;30m%%%%%%%%\033[0m\033[0;31m%%%%%%%%%%%%\033[0m\033[0;30m%%%%%%%%SSSS%%%%%%?\033[0m\033[0;32m????????????????????????????????????\033[0m\033[0;30m?%%%%SS\033[0m\033[0;37m+............\033[0m");
    $display("\033[0;37m...........*\033[0m\033[0;30m%%\033[0m\033[0;32m?????\033[0m\033[0;30m%%?\033[0m\033[0;32m??\033[0m\033[0;30m%%S%%\033[0m\033[0;31m?????????????????%%\033[0m\033[0;30m%%%%SSSSSSSS%%%%%%?\033[0m\033[0;32m???????????????????\033[0m\033[0;30m?%%%%%%%%%%\033[0m\033[0;31m%%%%??%%\033[0m\033[0;30m?\033[0m\033[0;37m............\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;32m?\033[0m\033[0;30m%%\033[0m\033[0;32m????\033[0m\033[0;30m?%%\033[0m\033[0;32m??\033[0m\033[0;30m%%S\033[0m\033[0;31m??????\033[0m\033[0;30mSSSSS%%\033[0m\033[0;31m%%%%?????????????%%\033[0m\033[0;30m%%SSSSSSSSSSSSSSSSSSSSSSSS%%%%\033[0m\033[0;31m%%??????%%\033[0m\033[0;30m%%\033[0m\033[0;37m;............\033[0m");
    $display("\033[0;37m...........;\033[0m\033[0;30m%%\033[0m\033[0;32m????\033[0m\033[0;30m%%%%\033[0m\033[0;32m??\033[0m\033[0;37m.\033[0m\033[0;31m???????????%%%%\033[0m\033[0;30m%%%%SSSSSSS%%%%\033[0m\033[0;31m%%%%?????????????????%%%%%%%%%%?????????????%%\033[0m\033[0;30m%%\033[0m\033[0;37m*,.............\033[0m");
    $display("\033[0;37m............\033[0m\033[0;32m*\033[0m\033[0;30m%%\033[0m\033[0;32m???\033[0m\033[0;30m%%%%\033[0m\033[0;32m??\033[0m\033[0;37m.\033[0m\033[0;30m%%\033[0m\033[0;31m?????????????????????%%%%%%\033[0m\033[0;30m%%SSSSSSSSSS%%%%\033[0m\033[0;31m%%%%???????????????%%%%\033[0m\033[0;30m%%SS#\033[0m\033[0;37m+,...............\033[0m");
    $display("\033[0;37m............,\033[0m\033[0;30m%%?\033[0m\033[0;32m??\033[0m\033[0;30m?\033[0m\033[0;32m???\033[0m\033[0;30m?S%%\033[0m\033[0;31m%%%%%%%%%%%%%%%%%%%%%%%%%%????????????????%%%%\033[0m\033[0;30m%%%%%%SSSSSSSSSSSSSSSSSSSSSS%%\033[0m\033[0;31m%%%%\033[0m\033[0;33m*\033[0m\033[0;37m................\033[0m");
    $display("\033[0;37m............,\033[0m\033[0;30mSS?\033[0m\033[0;32m???????\033[0m\033[0;30m%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;31m%%%%%%????????????????????????????????????%%?\033[0m\033[0;37m,...............\033[0m");
    $display("\033[0;37m............\033[0m\033[0;30m?S\033[0m\033[0;32m?\033[0m\033[0;30m%%%%\033[0m\033[0;32m?????????????????????????\033[0m\033[0;30m?%%%%SSSSSSS%%%%%%%%%%%%\033[0m\033[0;31m%%%%%%%%?????????????????%%%%?\033[0m\033[0;37m;,................\033[0m");
    $display("\033[0;37m...........*\033[0m\033[0;30m#%%\033[0m\033[0;32m??\033[0m\033[0;30m%%%%?\033[0m\033[0;32m???????????????????????????????\033[0m\033[0;30m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%SS%%\033[0m\033[0;31m???*\033[0m\033[0;33m*\033[0m\033[0;37m+;,...................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%\033[0m\033[0;30m%%%%\033[0m\033[0;32m??\033[0m\033[0;30m%%%%?\033[0m\033[0;32m?????????????????????????????????????????????\033[0m\033[0;30m?%%%%?\033[0m\033[0;37m*;,,,,........................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%\033[0m\033[0;30m%%%%%%%%%%%%\033[0m\033[0;32m???????????????????????????????????????\033[0m\033[0;30m%%%%%%?\033[0m\033[0;32m*\033[0m\033[0;37m+:...............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%\033[0m\033[0;30m%%%%SS%%%%\033[0m\033[0;32m??????????????????????????????\033[0m\033[0;30m?%%%%%%S%%\033[0m\033[0;36m*\033[0m\033[0;37m;,...................................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;30mSSSSS%%%%%%%%%%%%???????????\033[0m\033[0;32m???\033[0m\033[0;30m???\033[0m\033[0;32m?????\033[0m\033[0;30m??%%%%\033[0m\033[0;34m%%?\033[0m\033[0;37m+:..................................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%SS\033[0m\033[0;30mSSSSSSSSS%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;34m%%%%%%%%%%%%%%?\033[0m\033[0;37m+,...............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;36m*\033[0m\033[0;37m:.............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;37m;............................\033[0m");
    $display("\033[0;37m...........\033[0m\033[0;34m?%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%\033[0m\033[0;30mS\033[0m\033[0;37m+...........................\033[0m");
    $display("\033[0;37m...........::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::...........................\033[0m");
    $display("\033[0;37m....................................................................................................\033[0m");
    $display("\033[0;37m....................................................................................................\033[0m");
    $display("\033[31m \033[5m     //   / /     //   ) )     //   ) )     //   ) )     //   ) )\033[0m");
    $display("\033[31m \033[5m    //____       //___/ /     //___/ /     //   / /     //___/ /\033[0m");
    $display("\033[31m \033[5m   / ____       / ___ (      / ___ (      //   / /     / ___ (\033[0m");
    $display("\033[31m \033[5m  //           //   | |     //   | |     //   / /     //   | |\033[0m");
    $display("\033[31m \033[5m //____/ /    //    | |    //    | |    ((___/ /     //    | |\033[0m");

    /*$display("        ----------------------------               ");
    $display("        --                        --       |\__||  ");
    $display("        --  OOPS!!                --      / X,X  | ");
    $display("        --                        --    /_____   | ");
    $display("        --  \033[0;31mSimulation FAIL!!\033[m   --   /^ ^ ^ \\  |");
    $display("        --                        --  |^ ^ ^ ^ |w| ");
    $display("        ----------------------------   \\m___m__|_|");
    $display("\n");*/
end endtask

/*task display_pass; begin
        $display("\n");
        $display("\n");
        $display("        ----------------------------               ");
        $display("        --                        --       |\__||  ");
        $display("        --  Congratulations !!    --      / O.O  | ");
        $display("        --                        --    /_____   | ");
        $display("        --  \033[0;32mSimulation PASS!!\033[m     --   /^ ^ ^ \\  |");
        $display("        --                        --  |^ ^ ^ ^ |w| ");
        $display("        ----------------------------   \\m___m__|_|");
        $display("\n");
end endtask*/

task display_pass; begin
    $display("\033[0;37m......................................................,\033[0m\033[0;30m?%%%%%%\033[0m\033[0;37m+,.......................................\033[0m");
    $display("\033[0;37m.................................................,,::+\033[0m\033[0;30mS\033[0m\033[0;33m*::;?\033[0m\033[0;30m?\033[0m\033[0;33m*\033[0m\033[0;37m*+:...................................\033[0m");
    $display("\033[0;37m.........................................,+:...;\033[0m\033[0;30m?\033[0m\033[0;31m?\033[0m\033[0;33m*\033[0m\033[0;31m?\033[0m\033[0;30mSS\033[0m\033[0;33m+,,,::;+*\033[0m\033[0;31m?\033[0m\033[0;30mS\033[0m\033[0;37m*..................................\033[0m");
    $display("\033[0;37m........................................+\033[0m\033[0;30m%%\033[0m\033[0;37m.;.,*\033[0m\033[0;30m%%\033[0m\033[0;33m;,,,,,,,,,:;;:::;\033[0m\033[0;30m?\033[0m\033[0;37m*,................................\033[0m");
    $display("\033[0;37m.......................................;\033[0m\033[0;30mS\033[0m\033[0;33m:*\033[0m\033[0;30m%%??\033[0m\033[0;33m+,,:,,,,,;*+::;;;;;:*\033[0m\033[0;30m%%\033[0m\033[0;37m*,..............................\033[0m");
    $display("\033[0;37m.......................................+\033[0m\033[0;30m?\033[0m\033[0;33m,,,:,,;\033[0m\033[0;31m?*\033[0m\033[0;30m?\033[0m\033[0;33m*+*\033[0m\033[0;30m%%SS\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;33m+::::;;:;\033[0m\033[0;30m%%S\033[0m\033[0;37m:.............................\033[0m");
    $display("\033[0;37m.......................................:\033[0m\033[0;30mS\033[0m\033[0;33m:,,,:*\033[0m\033[0;30m?\033[0m\033[0;37m:,,;+;:,,:\033[0m\033[0;33m*\033[0m\033[0;30mS\033[0m\033[0;33m?+*\033[0m\033[0;30m?%%S%%\033[0m\033[0;33m;:\033[0m\033[0;31m?\033[0m\033[0;37m.:............................\033[0m");
    $display("\033[0;37m.......................................+.\033[0m\033[0;31m?\033[0m\033[0;33m;;+\033[0m\033[0;30m?\033[0m\033[0;37m*,,,,,,,,,,,,:\033[0m\033[0;33m+\033[0m\033[0;37m;;::;\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;33m;:\033[0m\033[0;30m%%S\033[0m\033[0;37m,...........................\033[0m");
    $display("\033[0;37m.......................................\033[0m\033[0;30mS\033[0m\033[0;33m+:\033[0m\033[0;30mS?\033[0m\033[0;37m*\033[0m\033[0;33m*\033[0m\033[0;37m:,,,,,,,,,;\033[0m\033[0;30m%%\033[0m\033[0;37m;,,,,,,,\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;33m;:+\033[0m\033[0;37m.;...........................\033[0m");
    $display("\033[0;37m.......................................+\033[0m\033[0;30m%%%%?\033[0m\033[0;37m,:,,,,,,,,,,,,;\033[0m\033[0;30m%%\033[0m\033[0;33m+\033[0m\033[0;37m,,,,;\033[0m\033[0;30mS%%\033[0m\033[0;33m;:;;\033[0m\033[0;37m.+...........................\033[0m");
    $display("\033[0;37m........................................\033[0m\033[0;30mSS\033[0m\033[0;37m,,,,,,,,,,,,,,,.,:,,,,+\033[0m\033[0;30m%%?\033[0m\033[0;33m+::+\033[0m\033[0;37m.;...........................\033[0m");
    $display("\033[0;37m.......................................:.:,:.\033[0m\033[0;30mS\033[0m\033[0;37m,,,,\033[0m\033[0;31m*\033[0m\033[0;37m,,,;\033[0m\033[0;30m?%%?\033[0m\033[0;37m:,,,,,;\033[0m\033[0;31m?\033[0m\033[0;30m??\033[0m\033[0;33m*:\033[0m\033[0;31m?\033[0m\033[0;37m.,...........................\033[0m");
    $display("\033[0;37m.......................................\033[0m\033[0;30m%%?\033[0m\033[0;37m,,:.\033[0m\033[0;30m%%\033[0m\033[0;37m,,,\033[0m\033[0;30m%%\033[0m\033[0;37m+,,,:;\033[0m\033[0;33m*\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m,,,,,;\033[0m\033[0;31m?\033[0m\033[0;30m?\033[0m\033[0;31m?\033[0m\033[0;30m?\033[0m\033[0;33m*\033[0m\033[0;37m.\033[0m\033[0;30m?\033[0m\033[0;37m............................\033[0m");
    $display("\033[0;37m.........,+\033[0m\033[0;33m*\033[0m\033[0;30m??%%\033[0m\033[0;37m:......................,.;,,,:,,:\033[0m\033[0;30mS\033[0m\033[0;37m*,,,,,,,,:,,,,,;\033[0m\033[0;33m**\033[0m\033[0;30m%%?\033[0m\033[0;37m..:............................\033[0m");
    $display("\033[0;37m........,\033[0m\033[0;30m?\033[0m\033[0;37m+:,,\033[0m\033[0;30m?%%\033[0m\033[0;37m......................:.:,,,,,:.\033[0m\033[0;30m%%\033[0m\033[0;37m.,,,,,,,,,,,,,,\033[0m\033[0;33m+*+\033[0m\033[0;37m+\033[0m\033[0;30mS\033[0m\033[0;37m.+.............................\033[0m");
    $display("\033[0;37m........\033[0m\033[0;33m*\033[0m\033[0;37m;,,,,\033[0m\033[0;30m?\033[0m\033[0;37m*......................:.:,,,,,,\033[0m\033[0;31m*\033[0m\033[0;37m.;,,,,,,,,,,,,,,:\033[0m\033[0;33m*\033[0m\033[0;37m,:.\033[0m\033[0;30mS\033[0m\033[0;37m..............................\033[0m");
    $display("\033[0;37m.......,\033[0m\033[0;30m?\033[0m\033[0;37m,,,,,\033[0m\033[0;30mS\033[0m\033[0;37m,......................:.;,,:,,,,::,,,,;\033[0m\033[0;30mS\033[0m\033[0;37m+,,,,,,,,,,,\033[0m\033[0;33m+\033[0m\033[0;37m.;.............................\033[0m");
    $display("\033[0;37m.......,\033[0m\033[0;30m%%\033[0m\033[0;37m,,,,;\033[0m\033[0;30m?\033[0m\033[0;37m.......................,.\033[0m\033[0;33m*\033[0m\033[0;37m,\033[0m\033[0;30mSS\033[0m\033[0;37m+;;::;;++*+\033[0m\033[0;34m*\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m:,,,,,,,,,\033[0m\033[0;33m+\033[0m\033[0;37m.;.............................\033[0m");
    $display("\033[0;37m........\033[0m\033[0;30m?\033[0m\033[0;37m;,,,:\033[0m\033[0;30m%%\033[0m\033[0;37m,.......................\033[0m\033[0;30m?\033[0m\033[0;37m.,\033[0m\033[0;30m?%%\033[0m\033[0;37m++;::::::;+*\033[0m\033[0;30m?S\033[0m\033[0;37m:,,,,,,:;\033[0m\033[0;33m*\033[0m\033[0;37m.*..............................\033[0m");
    $display("\033[0;37m......,,;.;,,,;\033[0m\033[0;30m?\033[0m\033[0;37m;,.....................:.\033[0m\033[0;30m?\033[0m\033[0;37m,::+\033[0m\033[0;30m???????\033[0m\033[0;37m*;,,;,,,,,:\033[0m\033[0;30m%%#?\033[0m\033[0;34m*\033[0m\033[0;37m:...............................\033[0m");
    $display("\033[0;37m...;\033[0m\033[0;30m?????S%%?\033[0m\033[0;33m*\033[0m\033[0;37m;,,\033[0m\033[0;33m+\033[0m\033[0;30m%%\033[0m\033[0;37m*,....................+.*.,,,+\033[0m\033[0;30m%%S\033[0m\033[0;37m+,,,,,,,,,,,;\033[0m\033[0;30mSS\033[0m\033[0;37m:..................................\033[0m");
    $display("\033[0;37m..;.;,,,,,,:;\033[0m\033[0;30m?%%\033[0m\033[0;33m+\033[0m\033[0;37m,:\033[0m\033[0;30mS%%\033[0m\033[0;37m,....................*.\033[0m\033[0;31m?\033[0m\033[0;37m,,,:;+:,,,,,,,,,:\033[0m\033[0;30m?\033[0m\033[0;37m.\033[0m\033[0;30mS\033[0m\033[0;37m;,..................................\033[0m");
    $display("\033[0;37m..*\033[0m\033[0;30mS\033[0m\033[0;37m.,,,,,,,,,:.;,:\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;30mS?\033[0m\033[0;37m+;:,............,,,+.\033[0m\033[0;30mS\033[0m\033[0;37m;,,,,,,,,,,,,:\033[0m\033[0;33m*\033[0m\033[0;30mS\033[0m\033[0;37m.\033[0m\033[0;33m*\033[0m\033[0;37m;\033[0m\033[0;33m+\033[0m\033[0;31m?\033[0m\033[0;30m%%\033[0m\033[0;37m+:,..............................\033[0m");
    $display("\033[0;37m..,\033[0m\033[0;30m?\033[0m\033[0;31m?\033[0m\033[0;37m+\033[0m\033[0;33m*\033[0m\033[0;31m?\033[0m\033[0;30m???\033[0m\033[0;33m*\033[0m\033[0;37m;::.\033[0m\033[0;33m*\033[0m\033[0;37m,,\033[0m\033[0;33m+\033[0m\033[0;37m.\033[0m\033[0;30m#\033[0m\033[0;34m?\033[0m\033[0;30m%%SS%%%%??\033[0m\033[0;34m*\033[0m\033[0;37m***\033[0m\033[0;34m*???\033[0m\033[0;30m???%%\033[0m\033[0;34m?\033[0m\033[0;30m%%S\033[0m\033[0;37m.\033[0m\033[0;30m%%\033[0m\033[0;37m+:,,,,,,,,,:;\033[0m\033[0;30m??\033[0m\033[0;37m,,,;.\033[0m\033[0;30m%%S%%\033[0m\033[0;37m*;,...........................\033[0m");
    $display("\033[0;37m...\033[0m\033[0;30m?%%\033[0m\033[0;37m;::::;+\033[0m\033[0;33m*\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;30m%%\033[0m\033[0;37m,,,\033[0m\033[0;33m*\033[0m\033[0;30mS%%\033[0m\033[0;36m+\033[0m\033[0;37m++++\033[0m\033[0;36m+********+++\033[0m\033[0;37m+++++\033[0m\033[0;30m%%\033[0m\033[0;31m?\033[0m\033[0;37m:+\033[0m\033[0;30m%%S?\033[0m\033[0;33m*+\033[0m\033[0;37m;:,,:\033[0m\033[0;33m+\033[0m\033[0;30m%%\033[0m\033[0;31m?\033[0m\033[0;37m,,,,\033[0m\033[0;30m%%#\033[0m\033[0;36m?\033[0m\033[0;34m??%%\033[0m\033[0;30mS%%\033[0m\033[0;37m*:.........................\033[0m");
    $display("\033[0;37m..,.;.,,,,...,:\033[0m\033[0;30m%%\033[0m\033[0;33m*\033[0m\033[0;37m,:\033[0m\033[0;30mS\033[0m\033[0;37m;\033[0m\033[0;33m*\033[0m\033[0;34m?\033[0m\033[0;37m+++++++++++++++++++++\033[0m\033[0;30m%%\033[0m\033[0;31m?\033[0m\033[0;37m,,:\033[0m\033[0;31m?\033[0m\033[0;37m...\033[0m\033[0;30mS%%%%%%%%\033[0m\033[0;31m?\033[0m\033[0;37m;,,,,\033[0m\033[0;30m%%\033[0m\033[0;37m.\033[0m\033[0;34m???????%%\033[0m\033[0;30mS%%\033[0m\033[0;37m;.......................\033[0m");
    $display("\033[0;37m...*\033[0m\033[0;30m%%\033[0m\033[0;37m++*\033[0m\033[0;33m**\033[0m\033[0;37m++;:,*\033[0m\033[0;30mS\033[0m\033[0;37m,\033[0m\033[0;33m*\033[0m\033[0;37m.,\033[0m\033[0;33m+\033[0m\033[0;34m%%\033[0m\033[0;36m?*+\033[0m\033[0;37m++++++++++++++++++\033[0m\033[0;36m*\033[0m\033[0;37m.;,,,:;\033[0m\033[0;33m+++\033[0m\033[0;37m;:,,,,,;\033[0m\033[0;30mS#\033[0m\033[0;34m??????????%%\033[0m\033[0;30mS%%\033[0m\033[0;37m;.....................\033[0m");
    $display("\033[0;37m....\033[0m\033[0;30m?S\033[0m\033[0;37m;;;;+\033[0m\033[0;33m*\033[0m\033[0;30m?%%S\033[0m\033[0;37m.;,\033[0m\033[0;33m+\033[0m\033[0;30m%%\033[0m\033[0;37m,\033[0m\033[0;33m*\033[0m\033[0;34m%%???\033[0m\033[0;36m**+\033[0m\033[0;37m++++++++++++++++\033[0m\033[0;36m*\033[0m\033[0;30m#\033[0m\033[0;33m+\033[0m\033[0;37m,,,,,,,,,,,:\033[0m\033[0;33m+\033[0m\033[0;30m%%#\033[0m\033[0;34m%%?????????????%%\033[0m\033[0;30m#%%\033[0m\033[0;37m:...................\033[0m");
    $display("\033[0;37m....\033[0m\033[0;30mS\033[0m\033[0;33m*\033[0m\033[0;37m.......,+.\033[0m\033[0;33m+\033[0m\033[0;37m,\033[0m\033[0;30m%%\033[0m\033[0;37m;:\033[0m\033[0;30mS\033[0m\033[0;34m???????\033[0m\033[0;36m***++++\033[0m\033[0;37m+\033[0m\033[0;34m?\033[0m\033[0;36m*\033[0m\033[0;37m+++++++\033[0m\033[0;30mS\033[0m\033[0;33m*\033[0m\033[0;37m,,,,,,,;\033[0m\033[0;33m*\033[0m\033[0;31m*\033[0m\033[0;30m%%SS\033[0m\033[0;34m%%?????????????????%%\033[0m\033[0;30mS\033[0m\033[0;37m*,.................\033[0m");
    $display("\033[0;37m....:\033[0m\033[0;30m#S\033[0m\033[0;31m*\033[0m\033[0;37m+;;;+*\033[0m\033[0;30m%%%%\033[0m\033[0;37m;\033[0m\033[0;30m?\033[0m\033[0;37m;;\033[0m\033[0;30m%%\033[0m\033[0;34m???????????????%%\033[0m\033[0;37m.\033[0m\033[0;34m?\033[0m\033[0;37m++++++\033[0m\033[0;36m+\033[0m\033[0;37m.;,,,,,,\033[0m\033[0;33m*\033[0m\033[0;30m#\033[0m\033[0;34m%%%%???????????????????????\033[0m\033[0;30mS%%\033[0m\033[0;37m:................\033[0m");
    $display("\033[0;37m.....,*\033[0m\033[0;30mS#%%%%??????\033[0m\033[0;33m+*\033[0m\033[0;30m%%\033[0m\033[0;34m????????%%%%%%\033[0m\033[0;30m%%%%%%\033[0m\033[0;34m?\033[0m\033[0;37m*+.\033[0m\033[0;34m?\033[0m\033[0;37m++++++\033[0m\033[0;34m?\033[0m\033[0;30mS\033[0m\033[0;37m,,,,,,,\033[0m\033[0;30mS\033[0m\033[0;34m%%\033[0m\033[0;36m?\033[0m\033[0;34m????????????????????????\033[0m\033[0;36m?\033[0m\033[0;34m%%\033[0m\033[0;30mS\033[0m\033[0;37m+...............\033[0m");
    $display("\033[0;37m........,:;++*\033[0m\033[0;30m??\033[0m\033[0;33m*\033[0m\033[0;30m%%S%%%%%%%%%%%%%%%%?\033[0m\033[0;36m*\033[0m\033[0;37m+;:,,..,.\033[0m\033[0;36m*\033[0m\033[0;37m++++++\033[0m\033[0;30m%%?\033[0m\033[0;37m,,,,,,:.\033[0m\033[0;34m?????????????????????????????\033[0m\033[0;30mS*\033[0m\033[0;37m..............\033[0m");
    $display("\033[0;37m...................,,,,,............,.\033[0m\033[0;34m?\033[0m\033[0;37m++++++\033[0m\033[0;30m#\033[0m\033[0;33m+\033[0m\033[0;37m,,,,,,;.\033[0m\033[0;34m??????????%%\033[0m\033[0;30mS\033[0m\033[0;34m%%?????????????????\033[0m\033[0;30mS%%\033[0m\033[0;37m,............\033[0m");
    $display("\033[0;37m....................................,.\033[0m\033[0;34m?\033[0m\033[0;37m++++++.;,,,,,,\033[0m\033[0;33m*\033[0m\033[0;30m#\033[0m\033[0;34m???????????\033[0m\033[0;30mSS#S%%\033[0m\033[0;34m???????????????\033[0m\033[0;30mS%%\033[0m\033[0;37m,...........\033[0m");
    $display("\033[0;32m \033[5m    //   ) )     // | |     //   ) )     //   ) )\033[m");
    $display("\033[0;32m \033[5m   //___/ /     //__| |    ((           ((\033[m");
    $display("\033[0;32m \033[5m  / ____ /     / ___  |      \\           \\\033[m");
    $display("\033[0;32m \033[5m //           //    | |        ) )          ) )\033[m");
    $display("\033[0;32m \033[5m//           //     | | ((___ / /    ((___ / /\033[m");
    $display("        ----------------------------               ");
    $display("        --                        --               ");
    $display("        --  Congratulations !!    --               ");
    $display("        --                        --               ");
    $display("        --  \033[0;32mSimulation PASS!!\033[m          ");
    $display("        --  total latency = %d        --               ",total_latency);
    $display("        --                        --               ");
    $display("        ----------------------------               ");
end endtask


endmodule